LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_Arith.ALL;
USE IEEE.STD_LOGIC_Unsigned.ALL;

ENTITY pipelining IS
PORT ( SWB       : IN   STD_LOGIC; 		--ģʽ����ֵ
       SWA	     : IN   STD_LOGIC;		--ģʽ����ֵ
	   SWC		 : IN   STD_LOGIC;		--Ϊ1ʱΪʵ��̨�����߼�ʵ��
	   clr       : IN   STD_LOGIC;		--��λ�źţ��͵�ƽ��Ч
       C	     : IN   STD_LOGIC;		--��λ��־ 
	   Z	     : IN   STD_LOGIC;		--���Ϊ���־
	   IRH	  	 : IN   STD_LOGIC_VECTOR(3 DOWNTO 0); --IR7,IR6,IR5,IR4��ָ�������
	   T3	 	 : IN   STD_LOGIC;		--T3ʱ��
	   W1	 	 : IN   STD_LOGIC;		--W1�������
	   W2	     : IN   STD_LOGIC;		--W2�������
	   W3   	 : IN   STD_LOGIC;		--W3�������
	   SELCTL	 : OUT   STD_LOGIC;		--Ϊ1ʱΪ����̨����
	   ABUS      : OUT   STD_LOGIC;		--Ϊ1ʱ�������������������
	   M         : OUT   STD_LOGIC;
	   S         : OUT   STD_LOGIC_VECTOR(3 DOWNTO 0); --S3,S2,S1,S0	   
	   SEL1      : OUT   STD_LOGIC; 	--SEL3��SEL2��SEL1��SEL0�൱�ڿ���̨��ʽʱ��ָ�������IR3��IR2��IR1��IR0
	   SEL0		 : OUT   STD_LOGIC;
	   SEL2		 : OUT   STD_LOGIC;
	   SEL3	     : OUT   STD_LOGIC;
	   DRW     	 : OUT   STD_LOGIC;		--Ϊ1ʱ������ۼ����͵�һ���ڶ��������Ĵ�������
	   SBUS      : OUT   STD_LOGIC;		--Ϊ1ʱ�������ݿ���ֵ����������
	   LIR       : OUT   STD_LOGIC;		--Ϊ1ʱ���Ӵ洢��������ָ����ָ��Ĵ���
	   MBUS      : OUT   STD_LOGIC;		--Ϊ1ʱ���Ӵ洢����������������������
	   MEMW      : OUT   STD_LOGIC;		--Ϊ1ʱ��T2д�洢����Ϊ0ʱ���洢��
	   LAR       : OUT   STD_LOGIC;		--Ϊ1ʱ��T2�������ؽ����������ϵĵ�ַ�����ַ�Ĵ���
	   ARINC     : OUT   STD_LOGIC;		--Ϊ1ʱ��T2�������ص�ַ�Ĵ�����1
	   LPC       : OUT   STD_LOGIC; 	--Ϊ1ʱ��T2�������ؽ����������ϵ����ݴ�����������PC
	   PCINC     : OUT   STD_LOGIC;		--Ϊ1ʱ��T2�������س����������1
	   PCADD	 : OUT	 STD_LOGIC;
	   CIN		 : OUT	 STD_LOGIC;
	   LONG		 : OUT   STD_LOGIC;
	   SHORT     : OUT   STD_LOGIC;
	   STOP		 : BUFFER STD_LOGIC;	--�۲�ʹ��
	   LDC		 : OUT   STD_LOGIC;		--Ϊ1ʱT3�������ر����λ
	   LDZ       : OUT   STD_LOGIC		--Ϊ1ʱT3�������ر�����Ϊ0��־	
	);
END pipelining;

ARCHITECTURE behavior OF pipelining IS 
SIGNAL ST0: STD_LOGIC;
SIGNAL SST0: STD_LOGIC;
SIGNAL SWCBA: STD_LOGIC_VECTOR(2 DOWNTO 0);
	

BEGIN
		
SWCBA <= SWC & SWB & SWA;
ST0_PROC: PROCESS(clr, T3)
	BEGIN
		IF clr = '0' THEN
			ST0 <= '0';
		ELSIF T3'EVENT AND T3 = '0' THEN
			IF SST0 = '1' THEN
				ST0 <= '1';
			END IF;
		END IF;
	END PROCESS;


OUT_SIG_PROC: PROCESS( SWCBA, IRH, W1, W2, W3, ST0, C, Z) 
  BEGIN
        --���ź�����Ĭ��ֵ
   SHORT 	<= '0';
   LONG		<= '0';
   CIN		<= '0';
   SELCTL   <= '0';
   ABUS     <= '0';
   SBUS	    <= '0';
   MBUS		<= '0';
   M        <= '0';
   S        <= "0000";
   SEL3		<= '0';
   SEL2		<= '0';
   SEL1     <= '0'; 
   SEL0		<= '0';
   DRW      <= '0';
   SBUS    <= '0';
   LIR      <= '0';
   MEMW     <= '0';
   	<='0';
   LAR      <= '0';
   ARINC    <= '0';
   LPC      <= '0';
   LDZ		<= '0';
   LDC		<= '0';
   STOP	    <= '0';
   PCINC	<= '0';
   SST0	<= '0';
   CASE SWCBA IS
		WHEN "000" =>   --ִ��ָ��
           CASE IRH IS  --ָ���
              
				WHEN "0000"=>
				LIR<=W1;
				PCINC<=W1;
				SHORT<=W1;

			  WHEN "0001" =>	--ADD
		   	LIR <= W1;  --ȡָ
        PCINC <= W1;
        SHORT<=W1;
				S <= "1001";
				CIN <= W1;
				ABUS <= W1;
				DRW <= W1;
				--LDC <= W1;
				LDZ <= W1;

				WHEN "0010" =>	--SUB
		   	LIR <= W1;  --ȡָ
        PCINC <= W1;
        SHORT<=W1;
				S <= "0110";
				ABUS <= W1;
				DRW <= W1;
				LDC <= W1;
				LDZ <= W1;

				WHEN "0011" =>	--AND
		   	LIR <= W1;  --ȡָ
        PCINC <= W1;
        SHORT<=W1;
				S <= "1011";
				M<=W1;
				ABUS <= W1;
				DRW <= W1;
				LDZ <= W1;
				
			  WHEN "0101" => --LD
				LAR <= W1;  --ȡָ
				M <= W1;
				S <= "1010";
				ABUS <= W1;
				LIR <= W2;
				PCINC<=W2;
				DRW <= W2;
				MBUS <= W2;
				
			  WHEN "0110" =>	--ST
				LAR <= W1;
				PCINC <= W2;
				M <= W2 OR W1;
				if W1 = '1' then
					S <= "1111";
				end if;
				if W2 = '1' then 
					S <= "1010";
				end if;
				ABUS <= W2 OR W1;
				LIR <= W2;
			    MEMW <= W2;
				
			  WHEN "0100" =>	--INC
				LIR <= W1;
				PCINC <= W1;
				SHORT<=W1;
				S <= "0000";
				ABUS <= W1;
				DRW <= W1;
				LDZ <= W1;
				LDC <= W1;
				
			  WHEN "1000" =>	--JZ
			    LIR <= ((NOT Z)AND W1) OR W2;
				PCINC <=  ((NOT Z)AND W1) OR W2;
				PCADD <= W1 AND Z;
				SHORT<=(NOT Z)AND W1;
				
			  WHEN "0111" =>	--JC
				LIR <= ((NOT C)AND W1) OR W2;  --ȡָ
		    PCINC <= ((NOT Z)AND W1) OR W2;
				PCADD <= W1 AND C;
				SHORT<=(NOT C)AND W1;
								
			  WHEN "1001" =>	--JMP
		   	    LIR <= W2;
				PCINC <= W2;
				LPC<=W1;
		        S <= "1111";
		        M <= W1;
		        ABUS <= W1;
				
			  WHEN "1110" =>	--STP
				STOP <= W1;
			
			  WHEN OTHERS =>--????????
				  LIR <= W1;
		      PCINC <= W1;
		          
					
		   END CASE;
		
		WHEN "001" =>	--д�洢��
		   SELCTL <= '1';
	  		SST0 <= NOT ST0 AND W1;
			SBUS <= W1;
	  		STOP <= W1;
			LAR  <= NOT ST0 AND W1;
			SHORT <= W1;
			MEMW <= ST0 AND W1;
			ARINC <= ST0 AND W1;
		   
			
		WHEN "010" =>	--���洢��
		   SBUS <= NOT ST0 AND W1;
		   LAR <= NOT ST0 AND W1;
		   STOP <= W1;
		   SST0 <= NOT ST0 AND W1;
		   SHORT <= W1 OR W2;
		   SELCTL <= '1';
		   MBUS <= ST0 AND W1;
		   ARINC <= W1 AND ST0;
		
		WHEN "011" =>	--���Ĵ���
		  SELCTL <= '1';
	  		STOP <= W1 OR W2;
			SEL3 <= W2;
			SEL2 <= W1 AND W2;
			SEL1<= W2;
			SEL0 <= W1 OR W2;
		  		 	
		WHEN "100" =>  --д�Ĵ���
			SELCTL	 <= '1';
	  		SST0 <= W2; 
			SBUS <= W1 OR W2;
	  		STOP <= W1 OR W2;
			DRW <= W1 OR W2;
			SEL3 <= (ST0 AND W1) OR (ST0 AND W2);
			SEL2 <= W2;
			SEL1<= (NOT ST0 AND	W1) OR (ST0 AND W2);
			SEL0 <= W1; 
		  
		WHEN OTHERS =>
			NULL;
	  END CASE;
		
	END PROCESS;
		
END behavior;